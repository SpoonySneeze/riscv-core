module alu (
    input [31:0] a, b,
    output [31:0] result
);
// Test comment for Git
//git test
endmodule